
 module decoder_7seg(
    input [3:0] hex_value,
    output reg [7:0] seg_7
    );
    
    always @(hex_value) begin
      case(hex_value) //숫자를 읽을 때는 underbar 유무 상관없다.
           4'b0000: seg_7 = 8'b0000_0011; //8'b11 //4'd3 //0
           4'b0001: seg_7 = 8'b1001_1111; //1
           4'b0010: seg_7 = 8'b0010_0101; //2
           4'b0011: seg_7 = 8'b0000_1101; //3
           4'b0100: seg_7 = 8'b1001_1001; //4
           4'b0101: seg_7 = 8'b0100_1001; //5
           4'b0110: seg_7 = 8'b0100_0001; //6
           4'b0111: seg_7 = 8'b0001_1011; //7
           4'b1000: seg_7 = 8'b0000_0001; //8
           4'b1001: seg_7 = 8'b0001_1001; //9
           4'b1010: seg_7 = 8'b0001_0001; //10,A
           4'b1011: seg_7 = 8'b1100_0001; //11,b
           4'b1100: seg_7 = 8'b0110_0011; //12,C
           4'b1101: seg_7 = 8'b1000_0101; //13,d
           4'b1110: seg_7 = 8'b0110_0001; //14,E
           4'b1111: seg_7 = 8'b0111_0001; //15,F      
       endcase
    end
       
 endmodule
